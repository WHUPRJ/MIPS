`include "defines.svh"

module instr_valid (
    input  word_t instr,
    output logic  valid
);

  always_comb
    casez (instr)
      32'b000000000000000000000?????001111: valid = 1'b1;  // SYNC (NOP)
      32'b00000000000???????????????000000: valid = 1'b1;  // SLL
      32'b00000000000???????????????000010: valid = 1'b1;  // SRL
      32'b00000000000???????????????000011: valid = 1'b1;  // SRA
      32'b000000???????????????00000000100: valid = 1'b1;  // SLLV
      32'b000000???????????????00000000110: valid = 1'b1;  // SRLV
      32'b000000???????????????00000000111: valid = 1'b1;  // SRAV
      32'b000000???????????????00000001010: valid = 1'b1;  // MOVZ
      32'b000000???????????????00000001011: valid = 1'b1;  // MOVN
      32'b000000?????000000000000000001000: valid = 1'b1;  // JR
      32'b000000?????00000?????00000001001: valid = 1'b1;  // JALR
      32'b000000????????????????????001100: valid = 1'b1;  // SYSCALL
      32'b000000????????????????????001101: valid = 1'b1;  // BREAK
      32'b0000000000000000?????00000010000: valid = 1'b1;  // MFHI
      32'b000000?????000000000000000010001: valid = 1'b1;  // MTHI
      32'b0000000000000000?????00000010010: valid = 1'b1;  // MFLO
      32'b000000?????000000000000000010011: valid = 1'b1;  // MTLO
      32'b000000??????????0000000000011000: valid = 1'b1;  // MULT
      32'b000000??????????0000000000011001: valid = 1'b1;  // MULTU
      32'b000000??????????0000000000011010: valid = 1'b1;  // DIV
      32'b000000??????????0000000000011011: valid = 1'b1;  // DIVU
      32'b000000???????????????00000100000: valid = 1'b1;  // ADD
      32'b000000???????????????00000100001: valid = 1'b1;  // ADDU
      32'b000000???????????????00000100010: valid = 1'b1;  // SUB
      32'b000000???????????????00000100011: valid = 1'b1;  // SUBU
      32'b000000???????????????00000100100: valid = 1'b1;  // AND
      32'b000000???????????????00000100101: valid = 1'b1;  // OR
      32'b000000???????????????00000100110: valid = 1'b1;  // XOR
      32'b000000???????????????00000100111: valid = 1'b1;  // NOR
      32'b000000???????????????00000101010: valid = 1'b1;  // SLT
      32'b000000???????????????00000101011: valid = 1'b1;  // SLTU
      32'b000000????????????????????110000: valid = 1'b1;  // TGE
      32'b000000????????????????????110001: valid = 1'b1;  // TGEU
      32'b000000????????????????????110010: valid = 1'b1;  // TLT
      32'b000000????????????????????110011: valid = 1'b1;  // TLTU
      32'b000000????????????????????110100: valid = 1'b1;  // TEQ
      32'b000000????????????????????110110: valid = 1'b1;  // TNE
      32'b000001?????00000????????????????: valid = 1'b1;  // BLTZ
      32'b000001?????00001????????????????: valid = 1'b1;  // BGEZ
      32'b000001?????01000????????????????: valid = 1'b1;  // TGEI
      32'b000001?????01001????????????????: valid = 1'b1;  // TGEIU
      32'b000001?????01010????????????????: valid = 1'b1;  // TLTI
      32'b000001?????01011????????????????: valid = 1'b1;  // TLTIU
      32'b000001?????01110????????????????: valid = 1'b1;  // TNEI
      32'b000001?????01100????????????????: valid = 1'b1;  // TEQI
      32'b000001?????10000????????????????: valid = 1'b1;  // BLTZAL
      32'b000001?????10001????????????????: valid = 1'b1;  // BGEZAL
      32'b000010??????????????????????????: valid = 1'b1;  // J
      32'b000011??????????????????????????: valid = 1'b1;  // JAL
      32'b000100??????????????????????????: valid = 1'b1;  // BEQ
      32'b000101??????????????????????????: valid = 1'b1;  // BNE
      32'b000110?????00000????????????????: valid = 1'b1;  // BLEZ
      32'b000111?????00000????????????????: valid = 1'b1;  // BGTZ
      32'b001000??????????????????????????: valid = 1'b1;  // ADDI
      32'b001001??????????????????????????: valid = 1'b1;  // ADDIU
      32'b001010??????????????????????????: valid = 1'b1;  // SLTI
      32'b001011??????????????????????????: valid = 1'b1;  // SLTIU
      32'b001100??????????????????????????: valid = 1'b1;  // ANDI
      32'b001101??????????????????????????: valid = 1'b1;  // ORI
      32'b001110??????????????????????????: valid = 1'b1;  // XORI
      32'b00111100000?????????????????????: valid = 1'b1;  // LUI
      32'b01000000000??????????00000000???: valid = 1'b1;  // MFC0
      32'b01000000100??????????00000000???: valid = 1'b1;  // MTC0
      32'b01000010000000000000000000000001: valid = 1'b1;  // TLBR
      32'b01000010000000000000000000000010: valid = 1'b1;  // TLBWI
      32'b01000010000000000000000000000110: valid = 1'b1;  // TLBWR
      32'b01000010000000000000000000001000: valid = 1'b1;  // TLBP
      32'b01000010000000000000000000011000: valid = 1'b1;  // ERET
      32'b011100??????????0000000000000000: valid = 1'b1;  // MADD
      32'b011100??????????0000000000000001: valid = 1'b1;  // MADDU
      32'b011100??????????0000000000000100: valid = 1'b1;  // MSUB
      32'b011100??????????0000000000000101: valid = 1'b1;  // MSUBU
      32'b011100???????????????00000000010: valid = 1'b1;  // MUL
      32'b100000??????????????????????????: valid = 1'b1;  // LB
      32'b100001??????????????????????????: valid = 1'b1;  // LH
      32'b100010??????????????????????????: valid = 1'b1;  // LWL
      32'b100011??????????????????????????: valid = 1'b1;  // LW
      32'b100100??????????????????????????: valid = 1'b1;  // LBU
      32'b100101??????????????????????????: valid = 1'b1;  // LHU
      32'b100110??????????????????????????: valid = 1'b1;  // LWR
      32'b101000??????????????????????????: valid = 1'b1;  // SB
      32'b101001??????????????????????????: valid = 1'b1;  // SH
      32'b101010??????????????????????????: valid = 1'b1;  // SWL
      32'b101011??????????????????????????: valid = 1'b1;  // SW
      32'b101110??????????????????????????: valid = 1'b1;  // SWR
      32'b101111?????00000????????????????: valid = 1'b1;  // I-Cache Index Invalid
      32'b101111?????01000????????????????: valid = 1'b1;  // I-Cache Index Store Tag
      32'b101111?????10000????????????????: valid = 1'b1;  // I-Cache Hit Invalid
      32'b101111?????00001????????????????: valid = 1'b1;  // D-Cache Index Writeback Invalid
      32'b101111?????01001????????????????: valid = 1'b1;  // D-Cache Index Store Tag
      32'b101111?????10001????????????????: valid = 1'b1;  // D-Cache Hit Invalid
      32'b101111?????10101????????????????: valid = 1'b1;  // D-Cache Hit Writeback Invalid
      32'b110011??????????????????????????: valid = 1'b1;  // PREF (NOP)
      default:                              valid = 1'b0;
    endcase
endmodule
